library verilog;
use verilog.vl_types.all;
entity led_text_tb is
end led_text_tb;
