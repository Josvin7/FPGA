library verilog;
use verilog.vl_types.all;
entity top_module_tb is
end top_module_tb;
